`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 03/24/2020 11:53:31 AM
// Design Name: 
// Module Name: tanh
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module tanh(
    input [4:0]count,
    output reg [31:0] partial
    );
//    reg [31:0]partial;
    always @(count)
    case(count)
        5'b00001: partial = 32'b00000000110010101110000000001101;
        5'b00010: partial = 32'b00000000010111100101010011100011;
        5'b00011: partial = 32'b00000000001011100110100010110010;
        5'b00100: partial = 32'b00000000000101110001110011111101;
        5'b00101: partial = 32'b00000000000010111000101110011010;
        5'b00110: partial = 32'b00000000000001011100010101110000;
        5'b00111: partial = 32'b00000000000000101110001010101100;
        5'b01000: partial = 32'b00000000000000010111000101010100;
        5'b01001: partial = 32'b00000000000000001011100010101010;
        5'b01010: partial = 32'b00000000000000000101110001010101;
        5'b01011: partial = 32'b00000000000000000010111000101010;
        5'b01100: partial = 32'b00000000000000000001011100010101;
        5'b01101: partial = 32'b00000000000000000000101110001010;
        5'b01110: partial = 32'b00000000000000000000010111000101;
        5'b01111: partial = 32'b00000000000000000000001011100010;
        5'b10000: partial = 32'b00000000000000000000000101110001;
        5'b10001: partial = 32'b00000000000000000000000010111000;
        5'b10010: partial = 32'b00000000000000000000000001011100;
        5'b10011: partial = 32'b00000000000000000000000000101110;
        5'b10100: partial = 32'b00000000000000000000000000010111;
        5'b10101: partial = 32'b00000000000000000000000000001011;
        5'b10110: partial = 32'b00000000000000000000000000000101;
        5'b10111: partial = 32'b00000000000000000000000000000010;
        5'b11000: partial = 32'b00000000000000000000000000000001;
        5'b11001: partial = 32'b00000000000000000000000000000000;
        5'b11010: partial = 32'b00000000000000000000000000000000;
        5'b11011: partial = 32'b00000000000000000000000000000000;
        5'b11100: partial = 32'b00000000000000000000000000000000;
        5'b11101: partial = 32'b00000000000000000000000000000000;
        5'b11110: partial = 32'b00000000000000000000000000000000;
    endcase
endmodule
